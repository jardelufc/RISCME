module imem(input  logic [31:0] a, output logic [31:0] rd);
  reg [31:0] ROM[255:0];
  initial begin
ROM[0]='hE04F000F;
ROM[1]='hE28020FF;
ROM[2]='hE5802804;
ROM[3]='hE5802804;
ROM[4]='hE5802804;
ROM[5]='hE5802804;
ROM[6]='hE5802804;
ROM[7]='hE28020FF;
ROM[8]='hE5802800;
ROM[9]='hE5802800;
ROM[10]='hE5802800;
ROM[11]='hE5802800;
ROM[12]='hE5802800;
ROM[13]='hE2802055;
ROM[14]='hE5802800;
ROM[15]='hE5802800;
ROM[16]='hE5802800;
ROM[17]='hE5802800;
ROM[18]='hE5802800;
ROM[19]='hE28020FF;
ROM[20]='hE5802800;
ROM[21]='hE5802800;
ROM[22]='hE5802800;
ROM[23]='hE5802800;
ROM[24]='hE5802800;
ROM[25]='hE2802055;
ROM[26]='hE5802800;
ROM[27]='hE5802800;
ROM[28]='hE5802800;
ROM[29]='hE5802800;
ROM[30]='hE5802800;
ROM[31]='hE28020FF;
ROM[32]='hE5802800;
ROM[33]='hE5802800;
ROM[34]='hE5802800;
ROM[35]='hE5802800;
ROM[36]='hE5802800;
ROM[37]='hE2802055;
ROM[38]='hE5802800;
ROM[39]='hE5802800;
ROM[40]='hE5802800;
ROM[41]='hE5802800;
ROM[42]='hE5802800;
ROM[43]='hE28020FF;
ROM[44]='hE5802800;
ROM[45]='hE5802800;
ROM[46]='hE5802800;
ROM[47]='hE5802800;
ROM[48]='hE5802800;
ROM[49]='hE2802055;
ROM[50]='hE5802800;
ROM[51]='hE5802800;
ROM[52]='hE5802800;
ROM[53]='hE5802800;
ROM[54]='hE5802800;
ROM[55]='hE28020FF;
ROM[56]='hE5802800;
ROM[57]='hE5802800;
ROM[58]='hE5802800;
ROM[59]='hE5802800;
ROM[60]='hE5802800;
ROM[61]='hE2802055;
ROM[62]='hE5802800;
ROM[63]='hE5802800;
ROM[64]='hE5802800;
ROM[65]='hE5802800;
ROM[66]='hE5802800;
ROM[67]='hE28020FF;
ROM[68]='hE5802800;
ROM[69]='hE5802800;
ROM[70]='hE5802800;
ROM[71]='hE5802800;
ROM[72]='hE5802800;
ROM[73]='hE2802055;
ROM[74]='hE5802800;
ROM[75]='hE5802800;
ROM[76]='hE5802800;
ROM[77]='hE5802800;
ROM[78]='hE58028;
  end
  assign rd = ROM[a[31:2]];
endmodule