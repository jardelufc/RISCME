ROM[0]='hE003E004;
ROM[1]='h00000031;
ROM[2]='h00000800;
ROM[3]='h1BF91BF8;
ROM[4]='h1BFC1BFB;
ROM[5]='h34AA3355;
ROM[6]='hD0F74323;
ROM[7]='h68436843;
ROM[8]='hE7F34798;
ROM[9]='hBF00BF00;
ROM[10]='hBF00BF00;
ROM[11]='hBF00BF00;
ROM[12]='h68811BF8;
ROM[13]='h1BFA6881;
ROM[14]='h600A32FF;
ROM[15]='h600A600A;
ROM[16]='h00004770;
